/*Copyright 2019-2021 T-Head Semiconductor Co., Ltd.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/
`define CLK_PERIOD          10
//`define JTLB_ENTRY_128
//`include "./cpu_cfig.h"
module cpu_mmu_mem_test_tb(
mmu_mem_passed
);
output mmu_mem_passed;
reg mmu_mem_passed;

//data array parameter

//==========================================================
//                  Parameter Definition
//==========================================================

//---------------------------------------------------------
// MMU Configuration
//---------------------------------------------------------
`define JTLB_ENTRY_1024
//`define JTLB_ENTRY_2048

`ifdef JTLB_ENTRY_1024
  `define JTLB_ADDR_WIDTH 8
`endif
`ifdef JTLB_ENTRY_2048
  `define JTLB_ADDR_WIDTH 9
`endif

`ifdef L1_CACHE_ECC
parameter LOCAL_DATA_DATA_WIDTH = 88;
parameter LOCAL_TAG_DATA_WIDTH  = 204;
`else
parameter LOCAL_DATA_DATA_WIDTH = 84;
parameter LOCAL_TAG_DATA_WIDTH  = 196;
`endif

//data
parameter LOCAL_DATA_ADDR_WIDTH  = `JTLB_ADDR_WIDTH;
parameter LOCAL_DATA_WE_WIDTH   = 4;
//tag
parameter LOCAL_TAG_ADDR_WIDTH = `JTLB_ADDR_WIDTH;
parameter LOCAL_TAG_WE_WIDTH   = 5;



//data array signal
reg [ LOCAL_DATA_ADDR_WIDTH-1 : 0 ] temp_data_addr_internal;
reg [ LOCAL_DATA_DATA_WIDTH-1 : 0 ] temp_data_din_internal ;
reg [ LOCAL_DATA_WE_WIDTH  -1 : 0 ] temp_data_wen_internal ;
reg                                 temp_data_cen0_internal ;
reg                                 temp_data_cen1_internal ;
reg                                 temp_data_CLK          ;
wire [ LOCAL_DATA_DATA_WIDTH-1 : 0] temp_data_q0_internal   ;
wire [ LOCAL_DATA_DATA_WIDTH-1 : 0] temp_data_q1_internal   ;
reg  [ LOCAL_DATA_DATA_WIDTH-1 : 0] golden_data      ;
reg  [ LOCAL_DATA_DATA_WIDTH-1 : 0] data0_mask   ;
reg  [ LOCAL_DATA_DATA_WIDTH-1 : 0] data0_mask_ff   ;
reg  [ LOCAL_DATA_DATA_WIDTH-1 : 0] data1_mask   ;

//tag array signal
reg [ LOCAL_TAG_ADDR_WIDTH-1 : 0 ] temp_tag_addr_internal;
reg [ LOCAL_TAG_DATA_WIDTH-1 : 0 ] temp_tag_din_internal ;
reg [ LOCAL_TAG_WE_WIDTH  -1 : 0 ] temp_tag_wen_internal ;
reg                                temp_tag_cen_internal ;
reg                                temp_tag_CLK          ;
wire [ LOCAL_TAG_DATA_WIDTH-1 : 0] temp_tag_q_internal   ;
reg  [ LOCAL_TAG_DATA_WIDTH-1 : 0] golden_tag      ;
reg  [ LOCAL_TAG_DATA_WIDTH-1 : 0] tag_mask   ;
reg  [ LOCAL_TAG_DATA_WIDTH-1 : 0] tag_mask_ff   ;

//gated cell clk
reg temp_forever_cpuclk      ;
reg temp_external_en         ;
reg temp_pad_yy_test_mode    ;
wire temp_xor_clk            ;


integer i;

initial 
begin
mmu_mem_passed = 1'b0;
//memory test
           temp_data_CLK               = 1'b0; 
           temp_data_cen0_internal     = 1'b1; 
           temp_data_cen1_internal     = 1'b0; 
           temp_data_wen_internal      = {LOCAL_DATA_WE_WIDTH{1'b1}};
           temp_data_addr_internal     = {LOCAL_DATA_ADDR_WIDTH{1'b0}};
           temp_data_din_internal      = {LOCAL_DATA_DATA_WIDTH{1'b0}};
           golden_data                 = {LOCAL_DATA_DATA_WIDTH{1'b0}};
           data0_mask                   = {LOCAL_DATA_DATA_WIDTH{1'b0}};
           #20
           @(posedge temp_data_CLK)

           //cen==1 test
           //$display("$$$$$$$$  data array  memory cen test cen ==1 test...                          $");   
           #0.1 temp_data_wen_internal   = {LOCAL_DATA_WE_WIDTH{1'b1}};
           #0.1 temp_data_cen0_internal  = 1'b1; 
           for(i=1;i<10;i=i+1)     //set address 1~9
           begin
               @(posedge temp_data_CLK)
                temp_data_addr_internal <= {LOCAL_DATA_ADDR_WIDTH{1'b0}} + i;
                temp_data_din_internal  <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + i;
                golden_data             <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + i;
           end

           @(posedge temp_data_CLK)

           //cen==1 test
           //$display("$$$$$$$$  data array  memory cen test cen ==1 test...                          $");   
           #0.1 temp_data_wen_internal   = {LOCAL_DATA_WE_WIDTH{1'b0}};
           #0.1 temp_data_cen0_internal  = 1'b1; 
           for(i=1;i<10;i=i+1)     //set address 1~9
           begin
               @(posedge temp_data_CLK)
                temp_data_addr_internal <= {LOCAL_DATA_ADDR_WIDTH{1'b0}} + i;
                temp_data_din_internal  <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + i;
                golden_data             <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + i;
               @(posedge temp_data_CLK)
               #0.1   
                   //$display("$address = %h temp_data_q0_internal = %h , golden_data =%h \n",temp_data_addr_internal,temp_data_q0_internal,golden_data);    
               if(temp_data_q0_internal !== golden_data)
               begin
                   //$display("$          Sorry, address %h memory write check fail ! @_@     $",temp_data_addr_internal);    
                   $finish;
               end
           end


           //cen==0 test
           //$display("$$$$$$$$$$  data array  memory cen test cen ==1  test passed                     $\n");   
           //$display("$$$$$$$$$$  data array  memory cen test  cen ==0 test...                         $");    
           #0.1 temp_data_wen_internal   = {LOCAL_DATA_WE_WIDTH{1'b1}};
           #0.1 temp_data_cen0_internal  = 1'b0; 

           for(i=10;i<15;i=i+1)     //set address 10 ~15
           begin
               @(posedge temp_data_CLK)
                temp_data_addr_internal <= {LOCAL_DATA_ADDR_WIDTH{1'b0}} + i;
                temp_data_din_internal  <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + i;
                golden_data             <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + i;
               @(posedge temp_data_CLK)
               #0.1   
                   //$display("$          address = %h temp_data_q0_internal = %h , golden_data =%h \n",temp_data_addr_internal,temp_data_q0_internal,golden_data);    
               if(temp_data_q0_internal === golden_data)
               begin
                   //$display("$          Sorry, address %h memory write check fail ! @_@     $",temp_data_addr_internal);    
                   $finish;
               end
           end


           //cen==1 test
           //$display("$$$$$$$$  data array  memory cen test cen ==1 test...                          $");   
           #0.1 temp_data_wen_internal   = {LOCAL_DATA_WE_WIDTH{1'b1}};
           #0.1 temp_data_cen1_internal  = 1'b1; 
           for(i=1;i<15;i=i+1)     //set address 1~9
           begin
               @(posedge temp_data_CLK)
                temp_data_addr_internal <= {LOCAL_DATA_ADDR_WIDTH{1'b0}} + i;
                temp_data_din_internal  <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + i;
                golden_data             <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + i;
           end

           #0.1 temp_data_wen_internal   = {LOCAL_DATA_WE_WIDTH{1'b0}};
           #0.1 temp_data_cen1_internal  = 1'b1; 
           for(i=1;i<15;i=i+1)     //set address 1~9
           begin
               @(posedge temp_data_CLK)
                temp_data_addr_internal <= {LOCAL_DATA_ADDR_WIDTH{1'b0}} + i;
                temp_data_din_internal  <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + i;
                golden_data             <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + i;
               @(posedge temp_data_CLK)
               #0.1   
                   //$display("$address = %h temp_data_q0_internal = %h , golden_data =%h \n",temp_data_addr_internal,temp_data_q0_internal,golden_data);    
               if(temp_data_q1_internal !== golden_data)
               begin
                   //$display("$          Sorry, address %h memory write check fail ! @_@     $",temp_data_addr_internal);    
                   $finish;
               end
           end


           //cen==0 test
           //$display("$$$$$$$$$$  data array  memory cen test cen ==1  test passed                     $\n");   
           //$display("$$$$$$$$$$  data array  memory cen test  cen ==0 test...                         $");    
           #0.1 temp_data_wen_internal   = {LOCAL_DATA_WE_WIDTH{1'b0}};
           #0.1 temp_data_cen1_internal  = 1'b1; 
           #0.1 temp_data_cen0_internal  = 1'b0; 

           for(i=10;i<15;i=i+1)     //set address 10 ~15
           begin
               @(posedge temp_data_CLK)
                temp_data_addr_internal <= {LOCAL_DATA_ADDR_WIDTH{1'b0}} + i;
                temp_data_din_internal  <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + i;
                golden_data             <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + i;
               @(posedge temp_data_CLK)
               #0.1   
                   //$display("$          address = %h temp_data_q0_internal = %h , golden_data =%h \n",temp_data_addr_internal,temp_data_q0_internal,golden_data);    
               if(temp_data_q1_internal !== golden_data)
               begin
                   //$display("$          Sorry, address %h memory write check fail ! @_@     $",temp_data_addr_internal);    
                   $finish;
               end
           end
          #0.1 temp_data_cen1_internal  = 1'b0; 

           //wen test
           //$display("$$$$$$$$$  data array  memory cen test  cen ==0 test passed                      $");    
           //$display("$$$$$$$$$  data array  memory wen test.......                                    $");    
           #0.1 temp_data_wen_internal   = {LOCAL_DATA_WE_WIDTH{1'b1}};
           #0.1 temp_data_cen0_internal   = 1'b1; 
          for(i=0;i<LOCAL_DATA_WE_WIDTH/2;i=i+1)
          begin
                 @(posedge temp_data_CLK)
                  temp_data_addr_internal <= {LOCAL_DATA_ADDR_WIDTH{1'b0}} ;
                  temp_data_wen_internal  <= {LOCAL_DATA_WE_WIDTH{1'b1}} <<i ; 
                  temp_data_din_internal  <= {20{1'b1}}<<56*i;
                  golden_data             <= {20{1'b1}}<<56*i;
                 @(posedge temp_data_CLK)
                 @(posedge temp_data_CLK)
                 #0.1 temp_data_wen_internal   <= {LOCAL_DATA_WE_WIDTH{1'b0}};
                       golden_data             <= temp_data_din_internal ;
                       data0_mask_ff           <= data0_mask;
                 @(posedge temp_data_CLK)
                  #0.1 
                    //  $display("$  address = %h temp_data_q0_internal = %h , golden_data =%h,wen=%h \n",temp_data_addr_internal,temp_data_q0_internal,(golden_data &(~data0_mask)),temp_data_wen_internal);    
                 if((temp_data_q0_internal & data0_mask_ff) !== (golden_data &(data0_mask_ff)) )
                 begin
                    //  $display("$  Sorry, temp_data_q0_internal = %h , golden_data =%h, wen=%h \n",temp_data_q0_internal,golden_data,temp_data_wen_internal);    
                      $finish;
                 end
           end
            
                      

          //write test
           //$display("$$$$$$$$$  data array  memory wen test passed                                    $");    
           //$display("$$$$$$$$$  data array  memory write test......                                   $");    
           @(posedge temp_data_CLK) //write address 0
           #0.1 temp_data_wen_internal   = {LOCAL_DATA_WE_WIDTH{1'b1}};
           #0.1 temp_data_cen0_internal   = 1'b1; 
           for(i=10;i<15;i = i+1)     //set address 10 ~15
           begin
           #0.1 temp_data_wen_internal   = {LOCAL_DATA_WE_WIDTH{1'b1}};
           #0.1 temp_data_cen0_internal   = 1'b1; 
               @(posedge temp_data_CLK)
                temp_data_addr_internal <= {LOCAL_DATA_ADDR_WIDTH{1'b0}} + i;
                temp_data_din_internal  <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + i;
                golden_data             <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + i;
               @(posedge temp_data_CLK)
               #0.1 temp_data_wen_internal   = {LOCAL_DATA_WE_WIDTH{1'b0}};
                    golden_data             <= temp_data_din_internal ;
               @(posedge temp_data_CLK)
               #0.1   
                   //$display("$          address = %h temp_data_q0_internal = %h , golden_data =%h \n",temp_data_addr_internal,temp_data_q0_internal,golden_data);    
               if(temp_data_q0_internal !== golden_data)
               begin
                   //$display("$          Sorry, address %h memory write check fail ! @_@     $",temp_data_addr_internal);    
                   $finish;
               end
           end

          //address width check
           //$display("$$$$$$$$  data array  memory read test passed                                    $");    
           //$display("$$$$$$$$  data array  memory address width test......                            $");    
           @(posedge temp_data_CLK) //write address 
           #0.1 temp_data_cen0_internal   = 1'b1; 
           @(posedge temp_data_CLK)
           temp_data_wen_internal  <= {LOCAL_DATA_WE_WIDTH{1'b1}};
           temp_data_addr_internal <= {LOCAL_DATA_ADDR_WIDTH{1'b0}} ;                // 0 address write bb
           temp_data_din_internal  <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + 8'hbb;
           golden_data             <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + 8'hbb;
           @(posedge temp_data_CLK)
           temp_data_wen_internal  <= {LOCAL_DATA_WE_WIDTH{1'b1}};
           temp_data_addr_internal <= { {1{1'b1}},{LOCAL_DATA_ADDR_WIDTH-1{1'b0}} } ; // 1/2 max address 
           temp_data_din_internal  <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + 8'haa;
           golden_data             <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + 8'haa;

           //read data in 1/2max address
           @(posedge temp_data_CLK)
           temp_data_wen_internal  <= {LOCAL_DATA_WE_WIDTH{1'b0}};
           temp_data_addr_internal <= { {1{1'b1}},{LOCAL_DATA_ADDR_WIDTH-1{1'b0}} } ; // 1/2 max address
           temp_data_din_internal  <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + 8'hff;
           golden_data             <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + 8'haa;
           @(posedge temp_data_CLK)
           #0.1   
           if(temp_data_q0_internal !== golden_data)
           begin
               //$display("$          Sorry, address %h memory read check fail ! @_@     $",temp_data_addr_internal);    
               $finish;
           end

           //read data in  address 0
           @(posedge temp_data_CLK)
           temp_data_wen_internal  <= {LOCAL_DATA_WE_WIDTH{1'b0}};
           temp_data_addr_internal <= {LOCAL_DATA_ADDR_WIDTH{1'b0}} ;                // 0 address write bb
           temp_data_din_internal  <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + 8'hff;
           golden_data             <= {LOCAL_DATA_DATA_WIDTH{1'b0}} + 8'hbb;
           @(posedge temp_data_CLK)
           #0.1   
           if(temp_data_q0_internal !== golden_data)
           begin
               //$display("$          Sorry, address %h memory read check fail ! @_@     $",temp_data_addr_internal);    
               $finish;
           end
           //$display("$$$$$$$$  data array  memory address width test passed                           $");    
           //$display("$$$$$$$$  data array  memory data width test......                               $");    
          //read data check
     
           @(posedge temp_data_CLK) //write address 
           #0.1 temp_data_cen0_internal   = 1'b1; 
           @(posedge temp_data_CLK)
           temp_data_wen_internal  <= {LOCAL_DATA_WE_WIDTH{1'b1}};
           temp_data_addr_internal <= {LOCAL_DATA_ADDR_WIDTH{1'b1}} ;
           temp_data_din_internal  <= {LOCAL_DATA_DATA_WIDTH{1'b1}} ;
           //golden_data             <= {LOCAL_DATA_DATA_WIDTH{1'b1}} ;
           @(posedge temp_data_CLK)
           #0.1 temp_data_wen_internal   = {LOCAL_DATA_WE_WIDTH{1'b0}};
                golden_data             <= temp_data_din_internal ;
           @(posedge temp_data_CLK)
           #0.1   
               //$display("$          address = %h temp_data_q0_internal = %h , golden_data =%h \n",temp_data_addr_internal,temp_data_q0_internal,golden_data);    
           if(temp_data_q0_internal !== golden_data)
           begin
               //$display("$          Sorry, address %h memory read check fail ! @_@     $",temp_data_addr_internal);    
               $finish;
           end
           //$display("$$$$$$$$  data array  memory data width test passed                          $");    
          //read data check
           //$display("$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$");
           //$display("$           data array test PASS!!!!!!!!!!!!!!!!!!!!                     $");    
           //$display("$           data array test PASS!!!!!!!!!!!!!!!!!!!!                     $");    
           //$display("$           data array test PASS!!!!!!!!!!!!!!!!!!!!                     $");    
           //$display("$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$");


           temp_tag_CLK               = 1'b0; 
           temp_tag_cen_internal      = 1'b0; 
           temp_tag_wen_internal      = {LOCAL_TAG_WE_WIDTH{1'b0}};
           temp_tag_addr_internal     = {LOCAL_TAG_ADDR_WIDTH{1'b0}};
           temp_tag_din_internal      = {LOCAL_TAG_DATA_WIDTH{1'b0}};
           golden_tag                 = {LOCAL_TAG_DATA_WIDTH{1'b0}};
           tag_mask                   = {LOCAL_TAG_DATA_WIDTH{1'b0}};

           #20
           @(posedge temp_tag_CLK)

           //cen==1 test
           //$display("$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$");
           //$display("$$$$$$$  tag array   memory cen test cen ==1 test...                  $");   
           //$display("$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$");
           #0.1 temp_tag_wen_internal   = {LOCAL_TAG_WE_WIDTH{1'b1}};
           #0.1 temp_tag_cen_internal  = 1'b1; 
           for(i=1;i<10;i=i+1)     //set address 1~9
           begin
           #0.1 temp_tag_wen_internal   = {LOCAL_TAG_WE_WIDTH{1'b1}};
           #0.1 temp_tag_cen_internal  = 1'b1; 
               @(posedge temp_tag_CLK)
                temp_tag_addr_internal <= {LOCAL_TAG_ADDR_WIDTH{1'b0}} + i;
                temp_tag_din_internal  <= {LOCAL_TAG_DATA_WIDTH{1'b0}} + i;
               // golden_tag             <= {LOCAL_TAG_DATA_WIDTH{1'b0}} + i;
               @(posedge temp_tag_CLK)
               #0.1 temp_tag_wen_internal   = {LOCAL_TAG_WE_WIDTH{1'b0}};
                    golden_tag             <= temp_tag_din_internal;
               @(posedge temp_tag_CLK)
               #0.1   
                   //$display("$address = %h temp_tag_q_internal = %h , golden_tag =%h \n",temp_tag_addr_internal,temp_tag_q_internal,golden_tag);    
               if(temp_tag_q_internal !== golden_tag)
               begin
                   //$display("$          Sorry, address %h memory write check fail ! @_@     $",temp_tag_addr_internal);    
                   $finish;
               end
           end


           //cen==0 test
           //$display("$$$$$$$$  tag array   memory cen test cen ==1  test passed                     $");   
           //$display("$$$$$$$$  tag array   memory cen test  cen ==0 test...                         $");    
           #0.1 temp_tag_wen_internal   = {LOCAL_TAG_WE_WIDTH{1'b0}};
           #0.1 temp_tag_cen_internal  = 1'b1; 

           for(i=10;i<15;i=i+1)     //set address 10 ~15
           begin
               @(posedge temp_tag_CLK)
                temp_tag_addr_internal <= {LOCAL_TAG_ADDR_WIDTH{1'b0}} + i;
                temp_tag_din_internal  <= {LOCAL_TAG_DATA_WIDTH{1'b0}} + i;
                golden_tag             <= {LOCAL_TAG_DATA_WIDTH{1'b0}} + i;
               @(posedge temp_tag_CLK)
               #0.1   
                   //$display("$          address = %h temp_tag_q_internal = %h , golden_tag =%h \n",temp_tag_addr_internal,temp_tag_q_internal,golden_tag);    
               if(temp_tag_q_internal === golden_tag)
               begin
                   //$display("$          Sorry, address %h memory write check fail ! @_@     $",temp_tag_addr_internal);    
                   $finish;
               end
           end



           //wen test
           //$display("$$$$$$$  tag array   memory cen test  cen ==0 test passed                      $");    
           //$display("$$$$$$$  tag array   memory wen test.......                                    $");    
           #0.1 temp_tag_wen_internal   = {LOCAL_TAG_WE_WIDTH{1'b1}};
           #0.1 temp_tag_cen_internal   = 1'b1; 
          for(i=0;i<LOCAL_TAG_WE_WIDTH + 1;i=i+1)
          begin
                 @(posedge temp_tag_CLK)
                  temp_tag_addr_internal <= {LOCAL_TAG_ADDR_WIDTH{1'b0}} ;
                  temp_tag_wen_internal  <= {LOCAL_TAG_WE_WIDTH{1'b1}} >>i ; 
                  temp_tag_din_internal  <= {LOCAL_TAG_DATA_WIDTH{1'b1}} ;
                 // golden_tag             <= {LOCAL_TAG_DATA_WIDTH{1'b1}} ;
                 @(posedge temp_tag_CLK)
                 @(posedge temp_tag_CLK)
                 #0.1 temp_tag_wen_internal  <= {LOCAL_TAG_WE_WIDTH{1'b0}};
                      golden_tag             <= temp_tag_din_internal;
                      tag_mask_ff            <= tag_mask;
                 @(posedge temp_tag_CLK)
                  #0.1 
                      //$display("$  address = %h temp_tag_q_internal = %h , golden_tag =%h,wen=%h \n",temp_tag_addr_internal,temp_tag_q_internal,(golden_tag &(tag_mask)),temp_tag_wen_internal);    
                 if((temp_tag_q_internal&tag_mask_ff) !== (golden_tag &(tag_mask_ff)) )
                 begin
                     // $display("$  temp_tag_q_internal = %h , golden_tag =%h, wen=%h (golden_tag &(~tag_mask)) =%h\n",temp_tag_q_internal,golden_tag,temp_tag_wen_internal, (golden_tag &(tag_mask)));    
                      $finish;
                 end
           end
            
                      

          //write test
           //$display("$$$$$$$$$  tag array   memory wen test passed                                    $");    
           //$display("$$$$$$$$$  tag array   memory write test......                                   $");    
           @(posedge temp_tag_CLK) //write address 0
           #0.1 temp_tag_wen_internal   = {LOCAL_TAG_WE_WIDTH{1'b1}};
           #0.1 temp_tag_cen_internal   = 1'b1; 
           for(i=10;i<15;i = i+1)     //set address 10 ~15
           begin
           #0.1 temp_tag_wen_internal   = {LOCAL_TAG_WE_WIDTH{1'b1}};
           #0.1 temp_tag_cen_internal   = 1'b1; 
               @(posedge temp_tag_CLK)
                temp_tag_addr_internal <= {LOCAL_TAG_ADDR_WIDTH{1'b0}} + i;
                temp_tag_din_internal  <= {LOCAL_TAG_DATA_WIDTH{1'b0}} + i;
                golden_tag             <= {LOCAL_TAG_DATA_WIDTH{1'b0}} + i;
               @(posedge temp_tag_CLK)
               #0.1 temp_tag_wen_internal   = {LOCAL_TAG_WE_WIDTH{1'b0}};
                    golden_tag             <= temp_tag_din_internal;
              @(posedge temp_tag_CLK)
               #0.1   
                   //$display("$          address = %h temp_tag_q_internal = %h , golden_tag =%h \n",temp_tag_addr_internal,temp_tag_q_internal,golden_tag);    
               if(temp_tag_q_internal !== golden_tag)
               begin
                   //$display("$          Sorry, address %h memory write check fail ! @_@     $",temp_tag_addr_internal);    
                   $finish;
               end
           end


          //address width check
           //$display("$$$$$$$$  tag array   memory read test passed                                    $");    
           //$display("$$$$$$$$  tag array   memory address width test......                            $");    
           @(posedge temp_tag_CLK) //write address 
           #0.1 temp_tag_cen_internal   = 1'b1; 
           //write address 0 
           @(posedge temp_tag_CLK)
           temp_tag_wen_internal  <= {LOCAL_TAG_WE_WIDTH{1'b1}};
           temp_tag_addr_internal <= {LOCAL_TAG_ADDR_WIDTH{1'b0}} ;
           temp_tag_din_internal  <= {LOCAL_TAG_DATA_WIDTH{1'b0}} + 8'hbb;
           golden_tag             <= {LOCAL_TAG_DATA_WIDTH{1'b0}} + 8'hbb;
           //write address 1/2 max address
           @(posedge temp_tag_CLK)
           temp_tag_wen_internal  <= {LOCAL_TAG_WE_WIDTH{1'b1}};
           temp_tag_addr_internal <= {{1'b1}, {LOCAL_TAG_ADDR_WIDTH-1{1'b0}} } ;
           temp_tag_din_internal  <= {LOCAL_TAG_DATA_WIDTH{1'b0}} + 8'haa;
           golden_tag             <= {LOCAL_TAG_DATA_WIDTH{1'b0}} + 8'haa;

           //read address 1/2 max address
           @(posedge temp_tag_CLK)
           temp_tag_wen_internal  <= {LOCAL_TAG_WE_WIDTH{1'b0}};
           temp_tag_addr_internal <= {{1'b1}, {LOCAL_TAG_ADDR_WIDTH-1{1'b0}} } ;
           temp_tag_din_internal  <= {LOCAL_TAG_DATA_WIDTH{1'b0}} + 8'hff;
           golden_tag             <= {LOCAL_TAG_DATA_WIDTH{1'b0}} + 8'haa;
           @(posedge temp_tag_CLK)
           #0.1   
           if(temp_tag_q_internal !== golden_tag)
           begin
               //$display("$          Sorry, address %h memory read check fail ! @_@     $",temp_tag_addr_internal);    
               $finish;
           end

           //read address 0
           @(posedge temp_tag_CLK)
           temp_tag_wen_internal  <= {LOCAL_TAG_WE_WIDTH{1'b0}};
           temp_tag_addr_internal <= {LOCAL_TAG_ADDR_WIDTH{1'b0}}  ;
           temp_tag_din_internal  <= {LOCAL_TAG_DATA_WIDTH{1'b0}} + 8'hff;
           golden_tag             <= {LOCAL_TAG_DATA_WIDTH{1'b0}} + 8'hbb;
           @(posedge temp_tag_CLK)
           #0.1   
           if(temp_tag_q_internal !== golden_tag)
           begin
               //$display("$          Sorry, address %h memory read check fail ! @_@     $",temp_tag_addr_internal);    
               $finish;
           end

           //$display("$$$$$$$  tag array   memory address width test passed                                $");    
           //$display("$$$$$$$  tag array   memory data width test......                                    $");    
          //read data check
     
           @(posedge temp_tag_CLK) //write address 
           #0.1 temp_tag_cen_internal   = 1'b1; 
           @(posedge temp_tag_CLK)
           temp_tag_wen_internal  <= {LOCAL_TAG_WE_WIDTH{1'b1}};
           temp_tag_addr_internal <= {LOCAL_TAG_ADDR_WIDTH{1'b1}} ;
           temp_tag_din_internal  <= {LOCAL_TAG_DATA_WIDTH{1'b1}} ;
           golden_tag             <= {LOCAL_TAG_DATA_WIDTH{1'b1}} ;
           @(posedge temp_tag_CLK)
           #0.1 temp_tag_wen_internal   = {LOCAL_TAG_WE_WIDTH{1'b0}};
                golden_tag             <= temp_tag_din_internal;
           @(posedge temp_tag_CLK)
           #0.1   
               //$display("$          address = %h temp_tag_q_internal = %h , golden_tag =%h \n",temp_tag_addr_internal,temp_tag_q_internal,golden_tag);    
           if(temp_tag_q_internal !== golden_tag)
           begin
               //$display("$          Sorry, address %h memory read check fail ! @_@     $",temp_tag_addr_internal);    
               $finish;
           end
           //$display("$$$$$$$  tag array   memory data width test passed                       $");    
          //read data check
           //$display("$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$");
           //$display("$           tag array test passed!!!!!!!!!!!!!!!!!!!!                    $");    
           //$display("$           tag array test passed!!!!!!!!!!!!!!!!!!!!                    $");    
           //$display("$           tag array test passed!!!!!!!!!!!!!!!!!!!!                    $");    
           //$display("$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$");

            #10
            mmu_mem_passed =1'b1;

end

////Dumping Control
//initial
//begin
//  $fsdbDumpfile("mmu_mem.fsdb");
//  $fsdbDumpon;
//  $fsdbDumpvars();
//  //$dumpfile("test.vcd");
//  //$dumpvars;
//end


always 
#(`CLK_PERIOD/2)  temp_data_CLK = ~temp_data_CLK;
always 
#(`CLK_PERIOD/2)  temp_tag_CLK = ~temp_tag_CLK;
//always 
//#(`CLK_PERIOD/2)  temp_dirty_CLK = ~temp_dirty_CLK;
always 
#(`CLK_PERIOD/2)  temp_forever_cpuclk = ~temp_forever_cpuclk;

always @(posedge temp_data_CLK)
begin
//data array mask
 data0_mask <= { {42{temp_data_wen_internal[1]}},{42{temp_data_wen_internal[0]}} };
 data1_mask <= { {42{temp_data_wen_internal[3]}},{42{temp_data_wen_internal[2]}} };
//tag array mask
tag_mask <= { {4{temp_tag_wen_internal[4]}} , {48{temp_tag_wen_internal[3]}},{48{temp_tag_wen_internal[2]}},{48{temp_tag_wen_internal[1]}} ,{48{temp_tag_wen_internal[0]}}};

end 



ct_mmu_jtlb_data_array x_px_mmu_da_smbist_wrap (
  .jtlb_data_idx               (  temp_data_addr_internal   ),
  .jtlb_data_cen0              (  temp_data_cen0_internal   ),
  .jtlb_data_cen1              (  temp_data_cen1_internal   ),
  .forever_cpuclk              (  temp_data_CLK             ),
  .jtlb_data_din               (  temp_data_din_internal    ),
  .jtlb_data_dout0             (  temp_data_q0_internal     ),
  .jtlb_data_dout1             (  temp_data_q1_internal     ),
  .jtlb_data_wen               (  temp_data_wen_internal    ),
  // .pad_yy_gate_clk_en_b          (  1'b0                      ),
  .pad_yy_icg_scan_en                 (   1'b1                     ),
  .cp0_mmu_icg_en            (  1'b1                      )
);

ct_mmu_jtlb_tag_array x_px_mmu_tag_smbist_wrap (
  .jtlb_tag_idx                    (temp_tag_addr_internal),
  .jtlb_tag_cen                    (temp_tag_cen_internal ),
  .forever_cpuclk                  (temp_tag_CLK          ),
  .jtlb_tag_din                    (temp_tag_din_internal ),
  .jtlb_tag_dout                   (temp_tag_q_internal   ),
  .jtlb_tag_wen                    (temp_tag_wen_internal ),
  // .pad_yy_gate_clk_en_b              (1'b0                  ),
  .pad_yy_icg_scan_en                 (   1'b1                     ),
  .cp0_mmu_icg_en                (1'b1                  )
);

endmodule
