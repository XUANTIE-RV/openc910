/*Copyright 2019-2021 T-Head Semiconductor Co., Ltd.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

// &ModuleBeg; @22
module ct_fadd_close_s0_d(
  close_adder0,
  close_adder1,
  close_eq,
  close_op_chg,
  close_sum_a_b,
  close_sum_b_a,
  ff1_pred,
  ff1_pred_onehot
);

// &Ports; @23
input   [52:0]  close_adder0;         
input   [52:0]  close_adder1;         
output          close_eq;             
output          close_op_chg;         
output  [52:0]  close_sum_a_b;        
output  [52:0]  close_sum_b_a;        
output  [5 :0]  ff1_pred;             
output  [52:0]  ff1_pred_onehot;      

// &Regs; @24
reg     [5 :0]  ff1_pred_50_0;        
reg     [52:0]  ff1_pred_onehot_50_0; 

// &Wires; @25
wire    [52:0]  close_adder0;         
wire    [52:0]  close_adder1;         
wire            close_eq;             
wire    [52:0]  close_ff1_a;          
wire    [52:0]  close_ff1_b;          
wire    [52:0]  close_ff1_c;          
wire    [52:0]  close_ff1_f;          
wire    [52:0]  close_ff1_g;          
wire    [52:0]  close_ff1_t;          
wire    [52:0]  close_ff1_z;          
wire            close_op_chg;         
wire    [53:0]  close_sum0;           
wire    [53:0]  close_sum1;           
wire    [52:0]  close_sum_a_b;        
wire    [52:0]  close_sum_b_a;        
wire    [5 :0]  ff1_pred;             
wire    [5 :0]  ff1_pred_52_51;       
wire    [5 :0]  ff1_pred_nz;          
wire    [52:0]  ff1_pred_nz_onehot;   
wire    [52:0]  ff1_pred_onehot;      
wire    [52:0]  ff1_pred_onehot_52_51; 

// &Force("nonport","close_sum1"); @26
// &Force("nonport","close_sum0"); @27
//close_sum0 for F0-F1
assign close_sum0[53:0]    = {1'b0,close_adder0[52:0]} 
                                       - {1'b0,close_adder1[52:0]};
assign close_sum1[53:0]    = {1'b0,close_adder1[52:0]} 
                                       - {1'b0,close_adder0[52:0]}; 
//notice that this situation, there is no need for m1, because the round
// m1 will never happen, there is no tail number used for rounding,
// here, it is different with the previous design


//close_sum select, keep sum not negative
//assign close_sum[52:0]     = (close_sum0[53])
//                           ? close_sum1[52:0]
//                           : close_sum0[52:0];
assign close_sum_a_b[52:0] = close_sum0[52:0];
assign close_sum_b_a[52:0] = close_sum1[52:0];
assign close_op_chg        = close_sum0[53];
assign close_eq            = !close_sum0[53] && !close_sum1[53];

//FF1 Logic of Close Path S0
//If predict first 1 set at r[n]
//Actual first 1 may set at r[n+1] or r[n]
//A and B are to oprand
assign close_ff1_a[52:0] = close_adder0[52:0];
assign close_ff1_b[52:0] = close_adder1[52:0];

//C = B && act_add || ~B && act_sub
assign close_ff1_c[52:0] = ~close_ff1_b[52:0];
//T = A^C  G=A&C  Z=(~A)&(~C)
assign close_ff1_t[52:0] = close_ff1_a[52:0] ^ close_ff1_c[52:0];
assign close_ff1_g[52:0] = close_ff1_a[52:0] & close_ff1_c[52:0];
assign close_ff1_z[52:0] = (~close_ff1_a[52:0]) & (~close_ff1_c[52:0]);
//F :
//fn-1 = En[gi(~zi-1) + zi(~gi-1)] + (~En)[gi(~gi-1) + zi(~zi-1)], En=act_sub
//f0   = t1(g0En+z0) + (~t1)(z0En+g0)
//fi   = ti+1[gi(~zi-1) + zi(~gi-1)] + (~ti+1)[gi(~gi-1) + zi(~zi-1)]
assign close_ff1_f[52]   =  ( close_ff1_g[52] & (~close_ff1_z[51])) | 
                            ( close_ff1_z[52] & (~close_ff1_g[51]));                          
assign close_ff1_f[0]    = (( close_ff1_t[1]) & (close_ff1_g[0] | close_ff1_z[0])) | 
                           ((~close_ff1_t[1]) & (close_ff1_z[0] | close_ff1_g[0]));
assign close_ff1_f[51:1] = (( close_ff1_t[52:2]) & ((close_ff1_g[51:1] & (~close_ff1_z[50:0])) | 
                            ( close_ff1_z[51:1]  & (~close_ff1_g[50:0]))))                     | 
                           ((~close_ff1_t[52:2]) & ((close_ff1_g[51:1] & (~close_ff1_g[50:0])) | 
                            ( close_ff1_z[51:1]  & (~close_ff1_z[50:0]))));                            

// &CombBeg; @73
always @( close_ff1_f[50:0])
begin
casez(close_ff1_f[50:0])
//  53'b1????_????????_????????_????????_????????_????????_???????? : 
//    ff1_pred_onehot_50_0[52:0] = 53'b10000_00000000_00000000_00000000_00000000_00000000_00000000;
//  53'b01???_????????_????????_????????_????????_????????_???????? : 
//    ff1_pred_onehot_50_0[52:0] = 53'b01000_00000000_00000000_00000000_00000000_00000000_00000000;
  51'b1??_????????_????????_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00100_00000000_00000000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd2;
  end
  51'b01?_????????_????????_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00010_00000000_00000000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd3;
  end
  51'b001_????????_????????_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00001_00000000_00000000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd4;
  end
  51'b000_1???????_????????_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_10000000_00000000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd5;
  end
  51'b000_01??????_????????_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_01000000_00000000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd6;
  end
  51'b000_001?????_????????_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00100000_00000000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd7;
  end
  51'b000_0001????_????????_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00010000_00000000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd8;
  end
  51'b000_00001???_????????_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00001000_00000000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd9;
  end
  51'b000_000001??_????????_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000100_00000000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd10;
  end
  51'b000_0000001?_????????_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000010_00000000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd11;
  end
  51'b000_00000001_????????_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000001_00000000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd12;
  end
  51'b000_00000000_1???????_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_10000000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd13;
  end
  51'b000_00000000_01??????_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_01000000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd14;
  end
  51'b000_00000000_001?????_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00100000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd15;
  end
  51'b000_00000000_0001????_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00010000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd16;
  end
  51'b000_00000000_00001???_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00001000_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd17;
  end
  51'b000_00000000_000001??_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000100_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd18;
  end
  51'b000_00000000_0000001?_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000010_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd19;
  end
  51'b000_00000000_00000001_????????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000001_00000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd20;
  end
  51'b000_00000000_00000000_1???????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_10000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd21;
  end
  51'b000_00000000_00000000_01??????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_01000000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd22;
  end
  51'b000_00000000_00000000_001?????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00100000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd23;
  end
  51'b000_00000000_00000000_0001????_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00010000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd24;
  end
  51'b000_00000000_00000000_00001???_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00001000_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd25;
  end
  51'b000_00000000_00000000_000001??_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000100_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd26;
  end
  51'b000_00000000_00000000_0000001?_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000010_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd27;
  end
  51'b000_00000000_00000000_00000001_????????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000001_00000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd28;
  end
  51'b000_00000000_00000000_00000000_1???????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_10000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd29;
  end
  51'b000_00000000_00000000_00000000_01??????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_01000000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd30;
  end
  51'b000_00000000_00000000_00000000_001?????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00100000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd31;
  end
  51'b000_00000000_00000000_00000000_0001????_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00010000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd32;
  end
  51'b000_00000000_00000000_00000000_00001???_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00001000_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd33;
  end
  51'b000_00000000_00000000_00000000_000001??_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000100_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd34;
  end
  51'b000_00000000_00000000_00000000_0000001?_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000010_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd35;
  end
  51'b000_00000000_00000000_00000000_00000001_????????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000001_00000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd36;
  end
  51'b000_00000000_00000000_00000000_00000000_1???????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_10000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd37;
  end
  51'b000_00000000_00000000_00000000_00000000_01??????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_01000000_00000000;
    ff1_pred_50_0[5:0]         = 6'd38;
  end
  51'b000_00000000_00000000_00000000_00000000_001?????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_00100000_00000000;
    ff1_pred_50_0[5:0]         = 6'd39;
  end
  51'b000_00000000_00000000_00000000_00000000_0001????_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_00010000_00000000;
    ff1_pred_50_0[5:0]         = 6'd40;
  end
  51'b000_00000000_00000000_00000000_00000000_00001???_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_00001000_00000000;
    ff1_pred_50_0[5:0]         = 6'd41;
  end
  51'b000_00000000_00000000_00000000_00000000_000001??_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_00000100_00000000;
    ff1_pred_50_0[5:0]         = 6'd42;
  end
  51'b000_00000000_00000000_00000000_00000000_0000001?_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_00000010_00000000;
    ff1_pred_50_0[5:0]         = 6'd43;
  end
  51'b000_00000000_00000000_00000000_00000000_00000001_???????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_00000001_00000000;
    ff1_pred_50_0[5:0]         = 6'd44;
  end
  51'b000_00000000_00000000_00000000_00000000_00000000_1??????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_00000000_10000000;
    ff1_pred_50_0[5:0]         = 6'd45;
  end
  51'b000_00000000_00000000_00000000_00000000_00000000_01?????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_00000000_01000000;
    ff1_pred_50_0[5:0]         = 6'd46;
  end
  51'b000_00000000_00000000_00000000_00000000_00000000_001????? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_00000000_00100000;
    ff1_pred_50_0[5:0]         = 6'd47;
  end
  51'b000_00000000_00000000_00000000_00000000_00000000_0001???? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_00000000_00010000;
    ff1_pred_50_0[5:0]         = 6'd48;
  end
  51'b000_00000000_00000000_00000000_00000000_00000000_00001??? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_00000000_00001000;
    ff1_pred_50_0[5:0]         = 6'd49;
  end
  51'b000_00000000_00000000_00000000_00000000_00000000_000001?? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_00000000_00000100;
    ff1_pred_50_0[5:0]         = 6'd50;
  end
  51'b000_00000000_00000000_00000000_00000000_00000000_0000001? : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_00000000_00000010;
    ff1_pred_50_0[5:0]         = 6'd51;
  end
  51'b000_00000000_00000000_00000000_00000000_00000000_00000001 : begin 
    ff1_pred_onehot_50_0[52:0] = 53'b00000_00000000_00000000_00000000_00000000_00000000_00000001;
    ff1_pred_50_0[5:0]         = 6'd52;
  end
  default : begin 
    ff1_pred_onehot_50_0[52:0] = {53{1'bx}};
    ff1_pred_50_0[5:0]         = {6{1'bx}};
  end
endcase
// &CombEnd; @288
end

assign ff1_pred_onehot_52_51[52:0] = (close_ff1_f[52])
                                   ? 53'b10000_00000000_00000000_00000000_00000000_00000000_00000000
                                   : 53'b01000_00000000_00000000_00000000_00000000_00000000_00000000;
assign ff1_pred_52_51[5:0]         = (close_ff1_f[52])
                                   ? 6'b0
                                   : 6'b1;

assign ff1_pred_nz_onehot[52:0] = (|close_ff1_f[52:51])
                                ? ff1_pred_onehot_52_51[52:0]
                                : ff1_pred_onehot_50_0[52:0];
assign ff1_pred_nz[5:0]         = (|close_ff1_f[52:51])
                                ? ff1_pred_52_51[5:0]
                                : ff1_pred_50_0[5:0];


assign ff1_pred_onehot[52:0] = ff1_pred_nz_onehot[52:0];
assign ff1_pred[5:0]         = ff1_pred_nz[5:0];
// &ModuleEnd; @307
endmodule


